// This is the unpowered netlist.
module cntr_example (wb_clk_i,
    wb_rst_i,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 output [37:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire clknet_0_wb_clk_i;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _047_ (.I(net1),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _048_ (.A1(net9),
    .A2(_020_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _049_ (.I(net1),
    .Z(_021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _050_ (.A1(net9),
    .A2(net10),
    .B(_021_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _051_ (.A1(net9),
    .A2(net10),
    .B(_022_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _052_ (.A1(net9),
    .A2(net10),
    .B(net11),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _053_ (.A1(net9),
    .A2(net10),
    .A3(net11),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _054_ (.A1(_021_),
    .A2(_024_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _055_ (.A1(_023_),
    .A2(_025_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _056_ (.A1(net12),
    .A2(_024_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _057_ (.A1(_020_),
    .A2(_026_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _058_ (.A1(net2),
    .A2(_020_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _059_ (.A1(net2),
    .A2(net13),
    .B(_021_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _060_ (.A1(net2),
    .A2(net13),
    .B(_027_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _061_ (.A1(net2),
    .A2(net13),
    .B(net14),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _062_ (.A1(net2),
    .A2(net13),
    .A3(net14),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _063_ (.A1(_021_),
    .A2(_029_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _064_ (.A1(_028_),
    .A2(_030_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _065_ (.A1(net15),
    .A2(_029_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _066_ (.A1(_020_),
    .A2(_031_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _067_ (.A1(net16),
    .A2(_020_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _068_ (.A1(net16),
    .A2(net17),
    .B(_021_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _069_ (.A1(net16),
    .A2(net17),
    .B(_032_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _070_ (.A1(net16),
    .A2(net17),
    .B(net18),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _071_ (.A1(net16),
    .A2(net17),
    .A3(net18),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _072_ (.A1(_021_),
    .A2(_034_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _073_ (.A1(_033_),
    .A2(_035_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _074_ (.A1(net19),
    .A2(_034_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _075_ (.A1(_020_),
    .A2(_036_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _076_ (.A1(net20),
    .A2(_020_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _077_ (.A1(net20),
    .A2(net21),
    .B(_021_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _078_ (.A1(net20),
    .A2(net21),
    .B(_037_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _079_ (.A1(net20),
    .A2(net21),
    .B(net3),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _080_ (.A1(net20),
    .A2(net21),
    .A3(net3),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _081_ (.A1(_021_),
    .A2(_039_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _082_ (.A1(_038_),
    .A2(_040_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _083_ (.A1(net4),
    .A2(_039_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _084_ (.A1(_020_),
    .A2(_041_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _085_ (.A1(net5),
    .A2(_020_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _086_ (.A1(net5),
    .A2(net6),
    .B(_021_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _087_ (.A1(net5),
    .A2(net6),
    .B(_042_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _088_ (.A1(net5),
    .A2(net6),
    .B(net7),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _089_ (.A1(net5),
    .A2(net6),
    .A3(net7),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _090_ (.A1(_021_),
    .A2(_044_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _091_ (.A1(_043_),
    .A2(_045_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _092_ (.A1(net8),
    .A2(_044_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _093_ (.A1(_020_),
    .A2(_046_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _094_ (.D(_000_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(net9));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _095_ (.D(_001_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(net10));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _096_ (.D(_002_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(net11));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _097_ (.D(_003_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(net12));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _098_ (.D(_004_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(net2));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _099_ (.D(_005_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(net13));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _100_ (.D(_006_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(net14));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _101_ (.D(_007_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(net15));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _102_ (.D(_008_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(net16));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _103_ (.D(_009_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(net17));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _104_ (.D(_010_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _105_ (.D(_011_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _106_ (.D(_012_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _107_ (.D(_013_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _108_ (.D(_014_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(net3));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _109_ (.D(_015_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(net4));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _110_ (.D(_016_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(net5));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _111_ (.D(_017_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(net6));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _112_ (.D(_018_),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(net7));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _113_ (.D(_019_),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(net8));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_23 (.ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_24 (.ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_25 (.ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_26 (.ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_27 (.ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_28 (.ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_29 (.ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_30 (.ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_31 (.ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_32 (.ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_33 (.ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_34 (.ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_35 (.ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_36 (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_523 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_524 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_525 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_526 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_527 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_528 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_529 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_530 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_531 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_532 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_533 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_534 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_535 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_536 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_537 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_538 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_539 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_540 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_541 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_542 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_543 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_544 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_545 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_546 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_547 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_548 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_549 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_550 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_551 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_552 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_553 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_554 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_555 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_556 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_557 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_558 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_559 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_560 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_561 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_562 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_563 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_564 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_565 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_566 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_567 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_568 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_569 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_570 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_571 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_572 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_573 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_574 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_575 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_576 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_577 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_578 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_579 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_580 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_581 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_582 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_583 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_584 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_585 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_586 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_587 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_588 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_589 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_590 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_591 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_592 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_593 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_594 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_595 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_596 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_597 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_598 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_599 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_600 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_601 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_602 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_603 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_604 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_605 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_606 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_607 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_608 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_609 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_610 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_611 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_612 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_613 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_614 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_615 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_616 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_617 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_618 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_619 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_620 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_621 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_622 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_623 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_624 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_625 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_626 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_627 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_628 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_629 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_630 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_631 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_632 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_633 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_634 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_635 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_636 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_637 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_638 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_639 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_640 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_641 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_642 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_643 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_644 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_645 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_646 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_647 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_648 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_649 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_650 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_651 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_652 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_653 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_654 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_655 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_656 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_657 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_658 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_659 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_660 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_661 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_662 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_663 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_664 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_665 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_666 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_667 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_668 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_669 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_670 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_671 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_672 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_673 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_674 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_675 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_676 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_677 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_678 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_679 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_680 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_681 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_682 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_683 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_684 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_685 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_686 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_687 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_688 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_689 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_690 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_691 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_692 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_693 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_694 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_695 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_696 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_697 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_698 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_699 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_700 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_701 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_702 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_703 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_704 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_705 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_706 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_707 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_708 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_709 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_710 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_711 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_712 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_713 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_714 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_715 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_716 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_717 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_718 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_719 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_720 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_721 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_722 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_723 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_724 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_725 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_726 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_727 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_728 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_729 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_730 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_731 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_732 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_733 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_734 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_735 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_736 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_737 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_738 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_739 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_740 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_741 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_742 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_743 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_744 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_745 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_746 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_7999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_8999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_9999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_10999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_11999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_12999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_13999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_14661 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(wb_rst_i),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output2 (.I(net2),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output3 (.I(net3),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output4 (.I(net4),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output5 (.I(net5),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output6 (.I(net6),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output7 (.I(net7),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output8 (.I(net8),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output9 (.I(net9),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output10 (.I(net10),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output11 (.I(net11),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output12 (.I(net12),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output13 (.I(net13),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output14 (.I(net14),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output15 (.I(net15),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output16 (.I(net16),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output17 (.I(net17),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output18 (.I(net18),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output19 (.I(net19),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output20 (.I(net20),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output21 (.I(net21),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel cntr_example_22 (.ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__094__D (.I(_000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__095__D (.I(_001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__096__D (.I(_002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__097__D (.I(_003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__098__D (.I(_004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__099__D (.I(_005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__100__D (.I(_006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__101__D (.I(_007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__102__D (.I(_008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__103__D (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__D (.I(_010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__105__D (.I(_011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__106__D (.I(_012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__107__D (.I(_013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__D (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__109__D (.I(_015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__110__D (.I(_016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__111__D (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__112__D (.I(_018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__113__D (.I(_019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__093__A1 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__085__A2 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__084__A1 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__076__A2 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__075__A1 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__067__A2 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__066__A1 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__058__A2 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__057__A1 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__048__A2 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__090__A1 (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__086__B (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__081__A1 (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__077__B (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__072__A1 (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__068__B (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__063__A1 (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__059__B (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__054__A1 (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__050__B (.I(_021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__051__B (.I(_022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__055__A1 (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__055__A2 (.I(_025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__057__A2 (.I(_026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__064__A1 (.I(_028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__065__A2 (.I(_029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__063__A2 (.I(_029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__064__A2 (.I(_030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__082__A1 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__083__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__081__A2 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__084__A2 (.I(_041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__091__A1 (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__092__A2 (.I(_044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__090__A2 (.I(_044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__091__A2 (.I(_045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__049__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__047__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output2_I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__062__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__061__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__060__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__059__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__058__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output3_I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__080__A3 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__079__B (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output4_I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__083__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output5_I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__089__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__088__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__087__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__086__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__085__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output6_I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__089__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__088__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__087__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__086__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output7_I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__089__A3 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__088__B (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output8_I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__092__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output9_I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__053__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__052__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__051__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__050__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__048__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output10_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__053__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__052__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__051__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__050__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output11_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__053__A3 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__052__B (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output12_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__056__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output13_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__062__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__061__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__060__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__059__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__062__A3 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__061__B (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__065__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__071__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__070__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__069__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__068__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__067__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__071__A2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__070__A2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__069__A2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__068__A2 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__071__A3 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__070__B (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__074__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__080__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__079__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__078__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__077__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__076__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__080__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__079__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__078__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__077__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__094__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__096__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__098__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__100__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__103__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__105__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__106__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__109__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__111__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__112__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__095__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__097__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__099__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__101__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__102__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__107__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__110__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__113__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_246_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_247_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_247_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_247_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_247_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_247_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_247_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_247_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_248_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_248_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_248_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_248_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_248_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_248_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_248_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_249_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_249_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_249_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_249_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_249_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_249_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_249_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_249_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_250_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_250_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_250_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_250_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_250_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_250_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_250_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_250_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_250_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_250_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_251_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_251_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_251_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_251_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_251_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_251_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_251_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_252_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_252_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_252_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_252_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_252_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_252_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_252_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_253_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_253_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_253_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_253_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_253_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_253_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_253_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_253_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_254_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_254_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_254_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_254_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_254_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_254_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_254_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_254_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_255_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_255_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_255_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_255_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_255_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_255_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_255_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_256_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_256_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_256_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_256_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_256_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_256_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_256_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_256_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_256_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_256_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_257_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_257_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_257_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_257_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_257_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_257_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_257_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_258_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_258_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_258_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_258_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_258_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_258_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_258_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_258_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_258_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_259_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_259_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_259_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_259_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_259_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_259_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_259_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_259_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_260_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_260_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_260_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_260_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_260_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_260_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_260_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_261_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_261_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_261_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_261_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_261_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_261_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_261_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_262_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_262_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_262_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_262_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_262_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_262_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_262_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_263_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_263_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_263_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_263_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_263_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_264_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_264_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_264_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_264_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_264_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_264_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_264_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_265_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_265_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_265_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_265_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_265_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_265_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_266_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_266_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_266_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_266_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_266_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_266_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_266_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_267_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_267_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_267_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_267_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_267_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_268_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_268_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_268_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_268_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_268_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_268_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_268_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_269_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_269_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_269_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_269_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_269_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_270_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_270_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_270_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_270_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_270_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_270_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_270_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_271_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_271_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_271_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_271_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_271_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_272_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_272_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_272_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_272_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_272_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_272_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_272_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_273_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_273_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_273_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_273_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_273_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_274_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_274_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_274_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_274_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_274_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_274_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_274_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_275_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_275_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_275_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_275_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_275_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_276_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_276_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_276_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_276_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_276_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_276_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_276_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_277_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_277_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_277_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_277_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_277_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_278_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_278_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_278_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_278_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_278_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_278_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_278_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_279_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_279_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_279_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_279_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_279_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_280_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_280_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_280_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_280_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_280_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_280_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_280_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_281_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_281_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_281_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_281_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_281_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_282_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_282_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_282_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_282_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_282_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_282_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_282_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_282_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_282_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_283_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_283_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_283_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_283_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_283_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_284_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_284_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_284_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_284_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_284_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_284_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_284_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_285_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_285_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_285_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_285_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_285_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_286_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_286_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_286_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_286_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_286_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_286_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_286_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_287_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_287_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_287_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_287_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_287_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_288_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_288_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_288_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_288_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_288_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_288_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_288_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_289_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_289_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_289_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_289_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_289_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_290_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_290_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_290_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_290_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_290_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_290_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_290_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_291_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_291_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_291_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_291_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_291_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_292_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_292_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_292_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_292_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_292_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_292_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_292_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_293_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_293_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_293_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_293_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_293_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_294_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_294_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_294_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_294_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_294_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_294_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_294_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_295_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_295_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_295_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_295_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_295_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_296_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_296_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_296_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_296_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_296_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_296_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_296_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_297_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_297_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_297_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_297_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_297_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_298_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_298_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_298_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_298_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_298_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_298_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_298_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_299_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_299_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_299_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_299_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_299_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_300_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_300_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_300_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_300_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_300_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_300_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_300_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_301_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_301_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_301_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_301_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_301_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_302_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_302_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_302_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_302_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_302_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_302_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_302_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_303_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_303_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_303_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_303_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_303_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_304_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_304_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_304_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_304_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_304_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_304_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_304_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_305_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_305_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_305_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_305_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_305_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_306_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_306_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_306_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_306_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_306_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_306_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_306_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_307_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_307_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_307_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_307_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_307_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_308_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_308_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_308_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_308_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_308_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_308_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_308_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_309_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_309_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_309_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_309_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_309_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_310_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_310_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_310_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_310_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_310_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_310_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_310_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_311_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_311_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_311_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_311_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_311_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_312_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_312_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_312_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_312_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_312_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_312_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_312_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_313_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_313_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_313_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_313_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_313_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_314_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_314_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_314_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_314_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_314_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_314_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_314_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_315_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_315_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_315_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_315_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_315_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_316_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_316_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_316_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_316_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_316_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_316_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_316_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_317_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_317_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_317_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_317_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_317_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_318_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_318_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_318_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_318_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_318_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_318_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_318_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_319_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_319_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_319_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_319_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_319_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_320_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_320_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_320_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_320_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_320_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_320_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_320_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_321_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_321_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_321_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_321_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_321_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_322_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_322_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_322_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_322_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_322_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_322_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_322_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_323_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_323_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_323_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_323_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_323_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_324_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_324_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_324_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_324_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_324_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_324_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_324_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_325_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_325_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_325_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_325_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_325_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_326_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_326_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_326_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_326_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_326_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_326_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_326_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_327_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_327_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_327_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_327_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_327_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_328_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_328_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_328_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_328_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_328_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_328_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_328_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_329_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_329_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_329_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_329_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_329_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_330_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_330_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_330_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_330_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_330_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_330_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_330_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_331_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_331_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_331_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_331_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_331_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_332_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_332_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_332_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_332_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_332_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_332_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_332_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_333_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_333_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_333_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_333_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_333_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_333_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_333_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_333_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_333_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_333_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_334_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_334_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_334_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_334_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_334_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_334_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_334_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_334_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_334_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_335_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_335_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_335_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_335_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_335_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_335_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_335_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_335_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_335_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_336_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_336_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_336_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_336_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_336_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_336_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_336_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_336_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_336_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_337_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_337_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_337_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_337_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_337_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_337_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_337_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_337_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_337_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_337_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_337_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_337_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_337_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_337_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_337_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_338_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_338_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_338_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_338_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_338_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_338_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_338_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_339_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_339_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_339_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_339_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_339_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_339_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_339_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_339_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_339_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_339_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_339_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_340_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_340_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_340_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_340_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_340_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_340_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_340_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_340_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_340_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_340_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_341_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_341_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_341_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_341_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_341_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_341_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_342_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_342_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_342_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_342_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_342_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_342_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_342_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_342_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_342_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_342_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_343_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_343_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_343_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_343_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_343_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_343_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_343_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_343_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_343_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_343_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_344_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_344_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_344_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_344_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_344_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_344_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_344_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_344_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_344_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_345_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_345_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_345_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_345_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_345_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_345_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_345_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_345_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_345_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_345_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_346_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_346_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_346_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_346_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_346_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_346_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_346_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_347_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_347_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_347_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_347_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_347_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_347_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_347_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_347_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_347_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_348_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_348_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_348_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_348_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_348_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_348_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_348_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_349_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_349_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_349_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_349_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_349_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_349_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_349_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_349_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_349_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_350_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_350_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_350_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_350_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_350_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_350_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_350_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_350_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_350_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_350_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_351_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_351_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_351_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_351_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_351_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_352_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_352_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_352_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_352_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_352_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_352_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_352_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_352_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_353_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_353_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_353_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_353_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_353_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_354_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_354_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_354_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_354_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_354_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_354_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_354_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_355_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_355_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_355_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_355_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_355_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_356_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_356_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_356_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_356_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_356_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_356_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_356_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_356_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_357_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_357_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_357_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_357_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_357_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_358_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_358_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_358_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_358_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_358_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_358_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_358_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_359_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_359_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_359_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_359_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_359_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_360_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_360_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_360_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_360_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_360_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_360_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_360_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_360_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_361_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_361_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_361_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_361_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_361_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_362_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_362_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_362_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_362_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_362_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_362_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_362_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_363_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_363_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_363_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_363_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_363_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_364_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_364_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_364_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_364_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_364_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_364_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_364_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_365_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_365_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_365_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_365_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_365_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_366_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_366_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_366_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_366_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_366_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_366_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_366_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_367_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_367_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_367_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_367_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_367_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_368_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_368_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_368_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_368_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_368_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_368_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_368_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_369_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_369_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_369_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_369_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_369_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_370_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_370_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_370_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_370_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_370_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_370_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_370_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_370_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_371_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_371_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_371_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_371_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_371_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_372_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_372_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_372_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_372_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_372_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_372_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_372_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_373_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_373_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_373_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_373_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_373_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_373_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_373_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_373_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_373_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_373_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_373_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_373_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_373_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_373_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_373_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_373_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_373_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_373_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_373_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_373_2651 ();
 assign io_out[20] = net22;
 assign io_out[21] = net23;
 assign io_out[22] = net24;
 assign io_out[23] = net25;
 assign io_out[24] = net26;
 assign io_out[25] = net27;
 assign io_out[26] = net28;
 assign io_out[27] = net29;
 assign io_out[28] = net30;
 assign io_out[29] = net31;
 assign io_out[30] = net32;
 assign io_out[31] = net33;
 assign io_out[32] = net34;
 assign io_out[33] = net35;
 assign io_out[34] = net36;
 assign io_out[35] = net37;
 assign io_out[36] = net38;
 assign io_out[37] = net39;
endmodule

